magic
tech sky130A
magscale 1 2
timestamp 1749490056
<< error_s >>
rect 19722 42861 19729 42891
rect 19756 42827 19763 42891
rect 18734 41090 18760 41110
rect 19447 29223 19454 29287
rect 19481 29257 19488 29287
rect 20478 27486 20504 27506
rect 7756 7188 7782 7208
rect 8744 5407 8751 5437
rect 8778 5407 8785 5471
<< mvpsubdiff >>
rect 3131 44155 3191 44189
rect 24839 44155 24899 44189
rect 3131 44129 3165 44155
rect 3131 31479 3165 31505
rect 24865 44129 24899 44155
rect 24865 31479 24899 31505
rect 3131 31445 3191 31479
rect 24839 31445 24899 31479
rect 2641 16985 2701 17019
rect 25029 16985 25089 17019
rect 2641 16959 2675 16985
rect 2641 4141 2675 4167
rect 25055 16959 25089 16985
rect 25055 4141 25089 4167
rect 2641 4107 2701 4141
rect 25029 4107 25089 4141
<< mvpsubdiffcont >>
rect 3191 44155 24839 44189
rect 3131 31505 3165 44129
rect 24865 31505 24899 44129
rect 3191 31445 24839 31479
rect 2701 16985 25029 17019
rect 2641 4167 2675 16959
rect 25055 4167 25089 16959
rect 2701 4107 25029 4141
<< locali >>
rect 3131 44155 3191 44189
rect 24839 44155 24899 44189
rect 3131 44129 24899 44155
rect 3165 44128 24865 44129
rect 3165 31526 3204 44128
rect 3244 44084 3296 44128
rect 24836 44084 24865 44128
rect 3244 44055 24865 44084
rect 3244 31571 3262 44055
rect 24773 44042 24865 44055
rect 24773 31571 24790 44042
rect 3244 31552 24790 31571
rect 3244 31526 3290 31552
rect 3165 31506 3290 31526
rect 24734 31510 24790 31552
rect 24834 31510 24865 44042
rect 24734 31506 24865 31510
rect 3165 31505 24865 31506
rect 3131 31479 24899 31505
rect 3131 31445 3191 31479
rect 24839 31445 24899 31479
rect 2641 16985 2701 17019
rect 25029 17018 25089 17019
rect 25029 16985 25095 17018
rect 2641 16959 25095 16985
rect 2675 16954 25055 16959
rect 2675 16916 2712 16954
rect 24926 16932 25055 16954
rect 24926 16916 24994 16932
rect 2675 16888 24994 16916
rect 2675 16864 2772 16888
rect 2675 4262 2700 16864
rect 2742 4262 2772 16864
rect 2675 4233 2772 4262
rect 24965 4254 24994 16888
rect 25038 4254 25055 16932
rect 24965 4233 25055 4254
rect 2675 4208 25055 4233
rect 2675 4168 2714 4208
rect 25024 4168 25055 4208
rect 2675 4167 25055 4168
rect 25089 4167 25095 16959
rect 2641 4141 25095 4167
rect 2641 4107 2701 4141
rect 25029 4107 25095 4141
rect 2643 4103 25095 4107
<< viali >>
rect 3204 31526 3244 44128
rect 3296 44084 24836 44128
rect 3290 31506 24734 31552
rect 24790 31510 24834 44042
rect 2712 16916 24926 16954
rect 2700 4262 2742 16864
rect 24994 4254 25038 16932
rect 2714 4168 25024 4208
<< metal1 >>
rect 3136 44181 3262 44186
rect 3136 44128 24899 44181
rect 3136 31914 3204 44128
rect 2305 31616 2311 31914
rect 2609 31616 3204 31914
rect 3136 31571 3204 31616
rect 3131 31526 3204 31571
rect 3244 44084 3296 44128
rect 24836 44084 24899 44128
rect 3244 44055 24899 44084
rect 3244 31571 3262 44055
rect 24773 44042 24899 44055
rect 24773 31571 24790 44042
rect 3244 31552 24790 31571
rect 3244 31526 3290 31552
rect 3131 31506 3290 31526
rect 24734 31510 24790 31552
rect 24834 31510 24899 44042
rect 24734 31506 24899 31510
rect 3131 31445 24899 31506
rect 2642 16954 25095 17018
rect 2642 16916 2712 16954
rect 24926 16932 25095 16954
rect 24926 16916 24994 16932
rect 2642 16888 24994 16916
rect 2642 16864 2772 16888
rect 2642 16484 2700 16864
rect 1976 16104 1982 16484
rect 2362 16104 2700 16484
rect 2642 4262 2700 16104
rect 2742 4262 2772 16864
rect 2642 4233 2772 4262
rect 24965 4254 24994 16888
rect 25038 4254 25095 16932
rect 24965 4233 25095 4254
rect 2642 4208 25095 4233
rect 2642 4168 2714 4208
rect 25024 4168 25095 4208
rect 2642 4108 25095 4168
rect 2643 4103 25095 4108
<< via1 >>
rect 2311 31616 2609 31914
rect 17576 43532 18276 43828
rect 20334 43536 21038 43862
rect 6330 42308 7044 42582
rect 8786 42426 9794 42582
rect 18162 29916 18888 30262
rect 20912 29922 21634 30246
rect 6176 28298 7152 28636
rect 8928 28284 9618 28622
rect 1982 16104 2362 16484
rect 17998 4918 18640 5188
rect 20456 4938 21408 5232
rect 6616 4466 7298 4760
rect 9372 4444 10060 4768
<< metal2 >>
rect 8300 44674 8356 44683
rect 8300 44609 8356 44618
rect 3068 44452 3128 44461
rect 2311 32517 2609 32526
rect 2311 31914 2609 32229
rect 2311 31610 2609 31616
rect 3068 31568 3128 44396
rect 7450 44270 7506 44279
rect 7450 44205 7506 44214
rect 6298 43152 7070 43172
rect 6298 42818 6316 43152
rect 7052 42818 7070 43152
rect 6298 42582 7070 42818
rect 7454 42628 7502 44205
rect 8304 42636 8352 44609
rect 12802 44538 12862 44547
rect 8744 43760 9822 43842
rect 8744 43486 8770 43760
rect 9794 43486 9822 43760
rect 8744 43126 9822 43486
rect 6298 42308 6330 42582
rect 7044 42308 7070 42582
rect 8744 42582 9824 43126
rect 8744 42426 8786 42582
rect 9794 42426 9824 42582
rect 8744 42394 9824 42426
rect 6298 42286 7070 42308
rect 12802 31568 12862 44482
rect 13544 44412 13604 44421
rect 13352 44146 13412 44155
rect 3064 31312 3128 31568
rect 7572 31534 7628 31543
rect 7572 31469 7628 31478
rect 12794 31534 12866 31568
rect 12794 31478 12796 31534
rect 12852 31478 12866 31534
rect 3064 31304 3124 31312
rect 3064 31248 3066 31304
rect 3122 31248 3124 31304
rect 3064 31246 3124 31248
rect 3066 31239 3122 31246
rect 6130 30640 7194 30708
rect 6130 30442 6152 30640
rect 7166 30442 7194 30640
rect 6130 28636 7194 30442
rect 7576 28648 7624 31469
rect 12794 31468 12866 31478
rect 8388 31304 8444 31313
rect 8388 31239 8444 31248
rect 8392 28636 8440 31239
rect 8890 31034 9670 31094
rect 8890 30858 8918 31034
rect 9654 30858 9670 31034
rect 6130 28298 6176 28636
rect 7152 28298 7194 28636
rect 6130 28266 7194 28298
rect 8890 28622 9670 30858
rect 13352 29538 13412 44090
rect 13544 31272 13604 44356
rect 18904 44274 18960 44283
rect 18904 44209 18960 44218
rect 19730 44270 19786 44279
rect 13760 44006 13820 44028
rect 13760 31452 13820 43950
rect 17538 43828 18652 43988
rect 17538 43532 17576 43828
rect 18276 43532 18652 43828
rect 18908 43788 18956 44209
rect 19730 44205 19786 44214
rect 19734 43778 19782 44205
rect 25396 44172 25456 44181
rect 20302 43862 21070 43976
rect 17538 43504 18652 43532
rect 18326 43166 18652 43504
rect 20302 43536 20334 43862
rect 21038 43762 21070 43862
rect 20302 43524 20336 43536
rect 21040 43524 21070 43762
rect 20302 43502 21070 43524
rect 18326 42828 18344 43166
rect 18634 42828 18652 43166
rect 18326 42806 18652 42828
rect 13760 31396 13762 31452
rect 13818 31396 13820 31452
rect 13760 31394 13820 31396
rect 20226 31452 20282 31461
rect 13762 31387 13818 31394
rect 20226 31387 20282 31396
rect 13544 31216 13546 31272
rect 13602 31216 13604 31272
rect 13544 31214 13604 31216
rect 19370 31272 19426 31281
rect 13546 31207 13602 31214
rect 19370 31207 19426 31216
rect 18144 30648 18916 31092
rect 18144 30440 18160 30648
rect 18898 30440 18916 30648
rect 18144 30262 18916 30440
rect 18144 29916 18162 30262
rect 18888 29916 18916 30262
rect 19374 30226 19422 31207
rect 20230 30164 20278 31387
rect 20892 31034 21664 31070
rect 20892 30860 20912 31034
rect 21644 30860 21664 31034
rect 20892 30246 21664 30860
rect 18144 29894 18916 29916
rect 20892 29922 20912 30246
rect 21634 29922 21664 30246
rect 20892 29898 21664 29922
rect 13352 29478 14054 29538
rect 8890 28284 8928 28622
rect 9618 28284 9670 28622
rect 8890 28256 9670 28284
rect 4446 17628 5564 17752
rect 4446 17320 4476 17628
rect 5546 17320 5564 17628
rect 4446 17254 5564 17320
rect 3991 17100 5985 17138
rect 3991 16768 4020 17100
rect 5966 16768 5985 17100
rect 3991 16668 5985 16768
rect 10241 17104 11142 17740
rect 10241 16776 10268 17104
rect 11118 16776 11142 17104
rect 10241 16750 11142 16776
rect 11516 17632 12656 17676
rect 11516 17306 11550 17632
rect 12630 17306 12656 17632
rect 11516 16664 12656 17306
rect 1982 16484 2362 16490
rect 1982 15920 2362 16104
rect 1982 15541 2362 15550
rect 6570 4760 7346 4794
rect 6570 4466 6616 4760
rect 7298 4466 7346 4760
rect 9324 4768 10094 4808
rect 3991 4222 5985 4434
rect 3991 3926 4014 4222
rect 5952 3926 5985 4222
rect 3991 3856 5985 3926
rect 6570 3442 7346 4466
rect 6570 3096 6600 3442
rect 7310 3096 7346 3442
rect 6570 3000 7346 3096
rect 7938 1934 7986 4488
rect 8784 3685 8832 4550
rect 9324 4444 9372 4768
rect 10060 4444 10094 4768
rect 8780 3676 8836 3685
rect 8780 3611 8836 3620
rect 9324 2694 10094 4444
rect 10662 3440 12656 4464
rect 13994 3676 14054 29478
rect 15576 17644 17570 18030
rect 15576 17298 15596 17644
rect 17554 17298 17570 17644
rect 15576 17254 17570 17298
rect 22247 17098 24241 18028
rect 25396 17580 25456 44116
rect 22247 16770 22258 17098
rect 24226 16770 24241 17098
rect 22247 16706 24241 16770
rect 24706 17520 25456 17580
rect 17928 5188 18696 5278
rect 16229 4206 17347 4922
rect 16229 3932 16264 4206
rect 17328 3932 17347 4206
rect 16229 3840 17347 3932
rect 17928 4918 17998 5188
rect 18640 4918 18696 5188
rect 20390 5232 21462 5298
rect 13994 3620 13996 3676
rect 14052 3620 14054 3676
rect 13994 3618 14054 3620
rect 13996 3611 14052 3618
rect 10662 3110 10702 3440
rect 12616 3110 12656 3440
rect 10662 3006 12656 3110
rect 17928 3444 18696 4918
rect 17928 3092 17954 3444
rect 18676 3092 18696 3444
rect 17928 3050 18696 3092
rect 9324 2410 9348 2694
rect 10068 2410 10094 2694
rect 9324 2340 10094 2410
rect 19084 2284 19132 4922
rect 19930 4051 19978 4954
rect 20390 4938 20456 5232
rect 21408 4938 21462 5232
rect 20390 4574 21462 4938
rect 19926 4042 19982 4051
rect 19926 3977 19982 3986
rect 20402 2696 21462 4574
rect 22024 3440 23142 4962
rect 24706 4042 24766 17520
rect 24706 3986 24708 4042
rect 24764 3986 24766 4042
rect 24706 3984 24766 3986
rect 24708 3977 24764 3984
rect 22024 3102 22054 3440
rect 23120 3102 23142 3440
rect 22024 3032 23142 3102
rect 20402 2404 20424 2696
rect 21434 2404 21462 2696
rect 20402 2326 21462 2404
rect 19084 2283 19332 2284
rect 19080 2274 19336 2283
rect 19080 2209 19336 2218
rect 7938 1933 8186 1934
rect 7934 1924 8190 1933
rect 7934 1859 8190 1868
<< via2 >>
rect 8300 44618 8356 44674
rect 3068 44396 3128 44452
rect 2311 32229 2609 32517
rect 7450 44214 7506 44270
rect 6316 42818 7052 43152
rect 12802 44482 12862 44538
rect 8770 43486 9794 43760
rect 4626 40842 5676 41726
rect 10440 39548 11460 40374
rect 13544 44356 13604 44412
rect 13352 44090 13412 44146
rect 7572 31478 7628 31534
rect 12796 31478 12852 31534
rect 3066 31248 3122 31304
rect 6152 30442 7166 30640
rect 8388 31248 8444 31304
rect 8918 30858 9654 31034
rect 18904 44218 18960 44274
rect 19730 44214 19786 44270
rect 13760 43950 13820 44006
rect 25396 44116 25456 44172
rect 20336 43536 21038 43762
rect 21038 43536 21040 43762
rect 20336 43524 21040 43536
rect 18344 42828 18634 43166
rect 15030 40862 16914 41722
rect 21690 39538 23584 40372
rect 13762 31396 13818 31452
rect 20226 31396 20282 31452
rect 13546 31216 13602 31272
rect 19370 31216 19426 31272
rect 18160 30440 18898 30648
rect 20912 30860 21644 31034
rect 4476 17320 5546 17628
rect 4020 16768 5966 17100
rect 10268 16776 11118 17104
rect 11550 17306 12630 17632
rect 1982 15550 2362 15920
rect 4014 3926 5952 4222
rect 6600 3096 7310 3442
rect 8780 3620 8836 3676
rect 15596 17298 17554 17644
rect 22258 16770 24226 17098
rect 16264 3932 17328 4206
rect 13996 3620 14052 3676
rect 10702 3110 12616 3440
rect 17954 3092 18676 3444
rect 9348 2410 10068 2694
rect 19926 3986 19982 4042
rect 24708 3986 24764 4042
rect 22054 3102 23120 3440
rect 20424 2404 21434 2696
rect 19080 2218 19336 2274
rect 7934 1868 8190 1924
<< metal3 >>
rect 8295 44676 8361 44679
rect 21770 44676 21776 44678
rect 8295 44674 21776 44676
rect 8295 44618 8300 44674
rect 8356 44618 21776 44674
rect 8295 44616 21776 44618
rect 8295 44613 8361 44616
rect 21770 44614 21776 44616
rect 21840 44614 21846 44678
rect 12797 44540 12867 44543
rect 22324 44540 22330 44542
rect 12797 44538 22330 44540
rect 12797 44482 12802 44538
rect 12862 44482 22330 44538
rect 12797 44480 22330 44482
rect 12797 44477 12867 44480
rect 22324 44478 22330 44480
rect 22394 44478 22400 44542
rect 3063 44454 3133 44457
rect 12400 44454 12406 44456
rect 3063 44452 12406 44454
rect 3063 44396 3068 44452
rect 3128 44396 12406 44452
rect 3063 44394 12406 44396
rect 3063 44391 3133 44394
rect 12400 44392 12406 44394
rect 12470 44392 12476 44456
rect 13539 44414 13609 44417
rect 22874 44414 22880 44416
rect 13539 44412 22880 44414
rect 13539 44356 13544 44412
rect 13604 44356 22880 44412
rect 13539 44354 22880 44356
rect 13539 44351 13609 44354
rect 22874 44352 22880 44354
rect 22944 44352 22950 44416
rect 7445 44272 7511 44275
rect 14594 44272 14600 44274
rect 7445 44270 14600 44272
rect 7445 44214 7450 44270
rect 7506 44214 14600 44270
rect 7445 44212 14600 44214
rect 7445 44209 7511 44212
rect 14594 44210 14600 44212
rect 14664 44210 14670 44274
rect 15140 44214 15146 44278
rect 15210 44276 15216 44278
rect 18899 44276 18965 44279
rect 15210 44274 18965 44276
rect 15210 44218 18904 44274
rect 18960 44218 18965 44274
rect 15210 44216 18965 44218
rect 15210 44214 15216 44216
rect 18899 44213 18965 44216
rect 19725 44272 19791 44275
rect 23420 44272 23426 44274
rect 19725 44270 23426 44272
rect 19725 44214 19730 44270
rect 19786 44214 23426 44270
rect 19725 44212 23426 44214
rect 19725 44209 19791 44212
rect 23420 44210 23426 44212
rect 23494 44210 23500 44274
rect 13347 44148 13417 44151
rect 23968 44148 23974 44150
rect 13347 44146 23974 44148
rect 13347 44090 13352 44146
rect 13412 44090 23974 44146
rect 13347 44088 23974 44090
rect 13347 44085 13417 44088
rect 23968 44086 23974 44088
rect 24038 44086 24044 44150
rect 24524 44112 24530 44176
rect 24594 44174 24600 44176
rect 25391 44174 25461 44177
rect 24594 44172 25461 44174
rect 24594 44116 25396 44172
rect 25456 44116 25461 44172
rect 24594 44114 25461 44116
rect 24594 44112 24600 44114
rect 25391 44111 25461 44114
rect 13755 44008 13825 44011
rect 15696 44008 15774 44010
rect 13755 44006 15774 44008
rect 13755 43950 13760 44006
rect 13820 44004 15774 44006
rect 13820 43950 15704 44004
rect 13755 43948 15704 43950
rect 13755 43945 13825 43948
rect 15696 43940 15704 43948
rect 15768 43940 15774 44004
rect 15696 43938 15774 43940
rect 218 43772 21115 43790
rect 218 43482 240 43772
rect 578 43762 21115 43772
rect 578 43760 20336 43762
rect 578 43486 8770 43760
rect 9794 43524 20336 43760
rect 21040 43524 21115 43762
rect 9794 43486 21115 43524
rect 578 43482 21115 43486
rect 218 43460 21115 43482
rect 782 43184 21178 43192
rect 782 43180 2678 43184
rect 782 42816 814 43180
rect 1188 42824 2678 43180
rect 2752 43166 21178 43184
rect 2752 43152 18344 43166
rect 2752 42824 6316 43152
rect 1188 42818 6316 42824
rect 7052 42828 18344 43152
rect 18634 42828 21178 43166
rect 7052 42818 21178 42828
rect 1188 42816 21178 42818
rect 782 42804 21178 42816
rect 1326 41740 23726 41768
rect 1326 40828 1424 41740
rect 1774 41726 23726 41740
rect 1774 40842 4626 41726
rect 5676 41722 23726 41726
rect 5676 40862 15030 41722
rect 16914 40862 23726 41722
rect 5676 40842 23726 40862
rect 1774 40828 23726 40842
rect 1326 40800 23726 40828
rect 794 40388 23826 40416
rect 794 39532 824 40388
rect 1170 40374 23826 40388
rect 1170 39548 10440 40374
rect 11460 40372 23826 40374
rect 11460 39548 21690 40372
rect 1170 39538 21690 39548
rect 23584 39538 23826 40372
rect 1170 39532 23826 39538
rect 794 39498 23826 39532
rect 783 32517 2614 32522
rect 783 32514 2311 32517
rect 783 32232 808 32514
rect 1188 32232 2311 32514
rect 783 32229 2311 32232
rect 2609 32229 2614 32517
rect 783 32224 2614 32229
rect 7567 31536 7633 31539
rect 12791 31536 12857 31539
rect 7567 31534 12857 31536
rect 7567 31478 7572 31534
rect 7628 31478 12796 31534
rect 12852 31478 12857 31534
rect 7567 31476 12857 31478
rect 7567 31473 7633 31476
rect 12791 31473 12857 31476
rect 13757 31454 13823 31457
rect 20221 31454 20287 31457
rect 13757 31452 20287 31454
rect 13757 31396 13762 31452
rect 13818 31396 20226 31452
rect 20282 31396 20287 31452
rect 13757 31394 20287 31396
rect 13757 31391 13823 31394
rect 20221 31391 20287 31394
rect 3061 31306 3127 31309
rect 8383 31306 8449 31309
rect 3061 31304 8449 31306
rect 3061 31248 3066 31304
rect 3122 31248 8388 31304
rect 8444 31248 8449 31304
rect 3061 31246 8449 31248
rect 3061 31243 3127 31246
rect 8383 31243 8449 31246
rect 13541 31274 13607 31277
rect 19365 31274 19431 31277
rect 13541 31272 19431 31274
rect 13541 31216 13546 31272
rect 13602 31216 19370 31272
rect 19426 31216 19431 31272
rect 13541 31214 19431 31216
rect 13541 31211 13607 31214
rect 19365 31211 19431 31214
rect 768 31042 21684 31054
rect 768 30846 814 31042
rect 1176 31034 21684 31042
rect 1176 30858 8918 31034
rect 9654 30860 20912 31034
rect 21644 30860 21684 31034
rect 9654 30858 21684 30860
rect 1176 30846 21684 30858
rect 768 30832 21684 30846
rect 200 30648 21694 30660
rect 200 30642 18160 30648
rect 200 30446 214 30642
rect 576 30640 18160 30642
rect 576 30446 6152 30640
rect 200 30442 6152 30446
rect 7166 30442 18160 30640
rect 200 30440 18160 30442
rect 18898 30440 21694 30648
rect 200 30424 21694 30440
rect 806 17650 24376 17660
rect 806 17294 822 17650
rect 1186 17644 24376 17650
rect 1186 17632 15596 17644
rect 1186 17628 11550 17632
rect 1186 17320 4476 17628
rect 5546 17320 11550 17628
rect 1186 17306 11550 17320
rect 12630 17306 15596 17632
rect 1186 17298 15596 17306
rect 17554 17298 24376 17644
rect 1186 17294 24376 17298
rect 806 17282 24376 17294
rect 1404 17114 24974 17124
rect 1404 16758 1420 17114
rect 1784 17104 24974 17114
rect 1784 17100 10268 17104
rect 1784 16768 4020 17100
rect 5966 16776 10268 17100
rect 11118 17098 24974 17104
rect 11118 16776 22258 17098
rect 5966 16770 22258 16776
rect 24226 16770 24974 17098
rect 5966 16768 24974 16770
rect 1784 16758 24974 16768
rect 1404 16746 24974 16758
rect 782 15920 2367 15925
rect 782 15904 1982 15920
rect 782 15568 820 15904
rect 1176 15568 1982 15904
rect 782 15550 1982 15568
rect 2362 15550 2367 15920
rect 782 15545 2367 15550
rect 1380 4232 17378 4250
rect 1380 3920 1428 4232
rect 1778 4222 17378 4232
rect 1778 3926 4014 4222
rect 5952 4206 17378 4222
rect 5952 3932 16264 4206
rect 17328 3932 17378 4206
rect 19921 4044 19987 4047
rect 24703 4044 24769 4047
rect 19921 4042 24769 4044
rect 19921 3986 19926 4042
rect 19982 3986 24708 4042
rect 24764 3986 24769 4042
rect 19921 3984 24769 3986
rect 19921 3981 19987 3984
rect 24703 3981 24769 3984
rect 5952 3926 17378 3932
rect 1778 3920 17378 3926
rect 1380 3890 17378 3920
rect 8775 3678 8841 3681
rect 13991 3678 14057 3681
rect 8775 3676 14057 3678
rect 8775 3620 8780 3676
rect 8836 3620 13996 3676
rect 14052 3620 14057 3676
rect 8775 3618 14057 3620
rect 8775 3615 8841 3618
rect 13991 3615 14057 3618
rect 790 3444 23265 3470
rect 790 3442 17954 3444
rect 790 3420 6600 3442
rect 790 3108 824 3420
rect 1174 3108 6600 3420
rect 790 3096 6600 3108
rect 7310 3440 17954 3442
rect 7310 3110 10702 3440
rect 12616 3110 17954 3440
rect 7310 3096 17954 3110
rect 790 3092 17954 3096
rect 18676 3440 23265 3444
rect 18676 3102 22054 3440
rect 23120 3102 23265 3440
rect 18676 3092 23265 3102
rect 790 3072 23265 3092
rect 218 2700 21488 2714
rect 218 2402 238 2700
rect 580 2696 21488 2700
rect 580 2694 20424 2696
rect 580 2410 9348 2694
rect 10068 2410 20424 2694
rect 580 2404 20424 2410
rect 21434 2404 21488 2696
rect 580 2402 21488 2404
rect 218 2384 21488 2402
rect 19075 2276 19341 2279
rect 27094 2276 27100 2278
rect 19075 2274 27100 2276
rect 19075 2218 19080 2274
rect 19336 2218 27100 2274
rect 19075 2216 27100 2218
rect 19075 2213 19341 2216
rect 27094 2214 27100 2216
rect 27364 2214 27370 2278
rect 7929 1926 8195 1929
rect 23214 1926 23220 1928
rect 7929 1924 23220 1926
rect 7929 1868 7934 1924
rect 8190 1868 23220 1924
rect 7929 1866 23220 1868
rect 7929 1863 8195 1866
rect 23214 1864 23220 1866
rect 23484 1864 23490 1928
<< via3 >>
rect 21776 44614 21840 44678
rect 22330 44478 22394 44542
rect 12406 44392 12470 44456
rect 22880 44352 22944 44416
rect 14600 44210 14664 44274
rect 15146 44214 15210 44278
rect 23426 44210 23494 44274
rect 23974 44086 24038 44150
rect 24530 44112 24594 44176
rect 15704 43940 15768 44004
rect 240 43482 578 43772
rect 814 42816 1188 43180
rect 2678 42824 2752 43184
rect 1424 40828 1774 41740
rect 824 39532 1170 40388
rect 808 32232 1188 32514
rect 814 30846 1176 31042
rect 214 30446 576 30642
rect 822 17294 1186 17650
rect 1420 16758 1784 17114
rect 820 15568 1176 15904
rect 1428 3920 1778 4232
rect 824 3108 1174 3420
rect 238 2402 580 2700
rect 27100 2214 27364 2278
rect 23220 1864 23484 1928
<< metal4 >>
rect 3006 44656 3066 45152
rect 3558 44656 3618 45152
rect 4110 44656 4170 45152
rect 4662 44656 4722 45152
rect 5214 44656 5274 45152
rect 5766 44656 5826 45152
rect 6318 44656 6378 45152
rect 6870 44656 6930 45152
rect 7422 44656 7482 45152
rect 7974 44656 8034 45152
rect 8526 44656 8586 45152
rect 9078 44656 9138 45152
rect 9630 44656 9690 45152
rect 10182 44656 10242 45152
rect 10734 44656 10794 45152
rect 11286 44656 11346 45152
rect 11838 44842 11898 45152
rect 12390 44842 12450 45152
rect 12942 44842 13002 45152
rect 13494 44842 13554 45152
rect 14046 45054 14106 45152
rect 14046 44952 14108 45054
rect 14598 45050 14658 45152
rect 15150 45106 15210 45152
rect 14598 44952 14662 45050
rect 11466 44750 13590 44842
rect 11466 44656 11558 44750
rect 2670 44564 11558 44656
rect 14048 44632 14108 44952
rect 12408 44572 14108 44632
rect 200 43772 600 44152
rect 200 43482 240 43772
rect 578 43482 600 43772
rect 200 30642 600 43482
rect 200 30446 214 30642
rect 576 30446 600 30642
rect 200 2700 600 30446
rect 200 2402 238 2700
rect 580 2402 600 2700
rect 200 1000 600 2402
rect 800 43180 1200 44152
rect 800 42816 814 43180
rect 1188 42816 1200 43180
rect 800 40388 1200 42816
rect 800 39532 824 40388
rect 1170 39532 1200 40388
rect 800 32514 1200 39532
rect 800 32232 808 32514
rect 1188 32232 1200 32514
rect 800 31042 1200 32232
rect 800 30846 814 31042
rect 1176 30846 1200 31042
rect 800 17650 1200 30846
rect 800 17294 822 17650
rect 1186 17294 1200 17650
rect 800 15904 1200 17294
rect 800 15568 820 15904
rect 1176 15568 1200 15904
rect 800 3420 1200 15568
rect 800 3108 824 3420
rect 1174 3108 1200 3420
rect 800 1000 1200 3108
rect 1400 41740 1800 44152
rect 2670 43184 2762 44564
rect 12408 44457 12468 44572
rect 12405 44456 12471 44457
rect 12405 44392 12406 44456
rect 12470 44392 12471 44456
rect 12405 44391 12471 44392
rect 14602 44275 14662 44952
rect 15148 44952 15210 45106
rect 15702 45006 15762 45152
rect 15702 44952 15766 45006
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 45022 21834 45152
rect 22326 45040 22386 45152
rect 21774 44952 21838 45022
rect 22326 44952 22392 45040
rect 22878 45032 22938 45152
rect 23430 45036 23490 45152
rect 22878 44952 22942 45032
rect 23430 44952 23492 45036
rect 23982 45030 24042 45152
rect 24534 45036 24594 45152
rect 15148 44279 15208 44952
rect 15145 44278 15211 44279
rect 14599 44274 14665 44275
rect 14599 44210 14600 44274
rect 14664 44210 14665 44274
rect 15145 44214 15146 44278
rect 15210 44214 15211 44278
rect 15145 44213 15211 44214
rect 14599 44209 14665 44210
rect 15706 44005 15766 44952
rect 21778 44679 21838 44952
rect 21775 44678 21841 44679
rect 21775 44614 21776 44678
rect 21840 44614 21841 44678
rect 21775 44613 21841 44614
rect 22332 44543 22392 44952
rect 22329 44542 22395 44543
rect 22329 44478 22330 44542
rect 22394 44478 22395 44542
rect 22329 44477 22395 44478
rect 22882 44417 22942 44952
rect 22879 44416 22945 44417
rect 22879 44352 22880 44416
rect 22944 44352 22945 44416
rect 22879 44351 22945 44352
rect 23432 44275 23492 44952
rect 23976 44952 24042 45030
rect 24532 44952 24594 45036
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 23425 44274 23495 44275
rect 23425 44210 23426 44274
rect 23494 44210 23495 44274
rect 23425 44209 23495 44210
rect 23976 44151 24036 44952
rect 24532 44177 24592 44952
rect 24529 44176 24595 44177
rect 23973 44150 24039 44151
rect 23973 44086 23974 44150
rect 24038 44086 24039 44150
rect 24529 44112 24530 44176
rect 24594 44112 24595 44176
rect 24529 44111 24595 44112
rect 23973 44085 24039 44086
rect 15703 44004 15769 44005
rect 15703 43940 15704 44004
rect 15768 43940 15769 44004
rect 15703 43939 15769 43940
rect 2670 42824 2678 43184
rect 2752 42824 2762 43184
rect 2670 42808 2762 42824
rect 1400 40828 1424 41740
rect 1774 40828 1800 41740
rect 1400 17114 1800 40828
rect 1400 16758 1420 17114
rect 1784 16758 1800 17114
rect 1400 4232 1800 16758
rect 1400 3920 1428 4232
rect 1778 3920 1800 4232
rect 1400 1000 1800 3920
rect 27099 2278 27365 2279
rect 27099 2214 27100 2278
rect 27364 2214 27365 2278
rect 27099 2213 27365 2214
rect 27102 2212 27362 2213
rect 23219 1928 23485 1929
rect 23219 1864 23220 1928
rect 23484 1864 23485 1928
rect 23219 1863 23485 1864
rect 23222 1862 23482 1863
rect 23422 200 23482 1862
rect 27302 200 27362 2212
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 200
use sky130_ef_ip__rc_osc_16M  sky130_ef_ip__rc_osc_16M_0 ../ip/sky130_ef_ip__rc_osc_16M/mag
timestamp 1749490056
transform 0 -1 13452 1 0 31680
box -24 680 10977 10082
use sky130_ef_ip__rc_osc_16M  sky130_ef_ip__rc_osc_16M_1
timestamp 1749490056
transform 0 1 2502 1 0 17748
box -24 680 10977 10082
use sky130_ef_ip__rc_osc_16M  sky130_ef_ip__rc_osc_16M_2
timestamp 1749490056
transform 0 -1 25086 -1 0 15801
box -24 680 10977 10082
use sky130_ef_ip__rc_osc_500k  sky130_ef_ip__rc_osc_500k_0 ../ip/sky130_ef_ip__rc_osc_500k/mag
timestamp 1749490056
transform 0 -1 24684 1 0 31634
box -24 -38 12264 10758
use sky130_ef_ip__rc_osc_500k  sky130_ef_ip__rc_osc_500k_1
timestamp 1749490056
transform 0 1 14526 1 0 18030
box -24 -38 12264 10758
use sky130_ef_ip__rc_osc_500k  sky130_ef_ip__rc_osc_500k_2
timestamp 1749490056
transform 0 -1 13706 -1 0 16664
box -24 -38 12264 10758
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1400 1000 1800 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
